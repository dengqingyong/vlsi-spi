`include "Internal_Ram.sv"
`include "packet.sv"
`include "master_host_if.sv"
`include "master_host_sequencer.sv"
`include "master_host_monitor.sv"
`include "master_host_driver.sv"
`include "master_host_agent.sv"
`include "master_host_env.sv"
`include "master_host_seq_lib.sv"

