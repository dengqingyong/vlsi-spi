class Internal_Ram;
	rand logic [7:0] ram [9:0];	//Internal RAM
endclass : Internal_Ram

