class Internal_Ram;
	rand logic [7:0] ram [1023:0];	//Internal RAM
endclass : Internal_Ram

